module sim();

wire [7:0] leds;
top top(.leds(leds));

endmodule