/*
This module provides FT245 synchronous FIFO functionality (e.g. for FT232H or FT2232H)
 */
 
 module ft245();
	 
endmodule
